
* Note: this is a placeholder for EPM
.SUBCKT EPM_Seq 2 3 4 5 6 7 8 9 10 11
* Forward (swap for reverse)
*A->B
*A->C
*A->D
*
*B->C
*B->D
*C->D
*                         0mS-10MS A->B ->C ->D                                              200ms-300ms B->C ->D A->D                          400-500ms B->A C->A D->A
VAP 3 2  PWL(000ms 0  10ms 5 10.00001ms 0  10.001001ms 5 10.002ms 5  10.002001ms 0  20.00000ms 0  20.000001ms 5 20.002ms 5  20.002001ms 0   30.000001ms 0  30.001001ms 0 30.002ms 0  30.002001ms 0   )
VAN 4 2  PWL(000ms 0  10ms 0 10.00001ms 0  10.001001ms 0 10.002ms 0  10.002001ms 0  20.00000ms 0  20.000001ms 0 20.002ms 0  20.002001ms 0   30.000001ms 0  30.001001ms 5 30.002ms 5  30.002001ms 0   )
VBP 5 2  PWL(000ms 0  10ms 0 10.00001ms 0  10.001001ms 0 10.002ms 0  10.002001ms 0  20.00000ms 0  20.000001ms 5 20.002ms 5  20.002001ms 0   30.000001ms 0  30.001001ms 5 30.002ms 5  30.002001ms 0   )
VBN 6 2  PWL(000ms 0  10ms 5 10.00001ms 0  10.001001ms 5 10.002ms 5  10.002001ms 0  20.00000ms 0  20.000001ms 0 20.002ms 0  20.002001ms 0   30.000001ms 0  30.001001ms 0 30.002ms 0  30.002001ms 0   )
VCP 7 2  PWL(000ms 0  10ms 0 10.00001ms 0  10.001001ms 0 10.002ms 0  10.002001ms 0  20.00000ms 0  20.000001ms 0 20.002ms 0  20.002001ms 0   30.000001ms 0  30.001001ms 5 30.002ms 5  30.002001ms 0   )
VCN 8 2  PWL(000ms 0  10ms 5 10.00001ms 0  10.001001ms 5 10.002ms 5  10.002001ms 0  20.00000ms 0  20.000001ms 5 20.002ms 5  20.002001ms 0   30.000001ms 0  30.001001ms 0 30.002ms 0  30.002001ms 0    )
VDP 9 2  PWL(000ms 0  10ms 0 10.00001ms 0  10.001001ms 0 10.002ms 0  10.002001ms 0  20.00000ms 0  20.000001ms 0 20.002ms 0  20.002001ms 0   30.000001ms 0  30.001001ms 5 30.002ms 5  30.002001ms 0    )
VDN 10 2 PWL(000ms 0  10ms 5 10.00001ms 0  10.001001ms 5 10.002ms 5  10.002001ms 0  20.00000ms 0  20.000001ms 5 20.002ms 5  20.002001ms 0   30.000001ms 0  30.001001ms 0 30.002ms 0  30.002001ms 0   )

VEnable 11 2 5V
*VBP 6 2  PWL(000ms 5  200ms 5 200.001ms 0  400ms 0 400.001ms 5   600ms 5 600.001ms 0  800ms 0 800.001ms 5  1000ms 5 1000.001ms 0  1200ms 0 1200.001ms 5)
*VBN 4 2  PWL(000ms 0  200ms 0 200.001ms 5  400ms 5 400.001ms 0   600ms 0 600.001ms 5  800ms 5 800.001ms 0  1000ms 0 1000.001ms 5  1200ms 5 1200.001ms 0)

.ENDS EPM_Seq
