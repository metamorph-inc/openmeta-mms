* L_LINEAR
* SPICE model of a linear inductor.
*
*
*----------------------------------------------
*  External Pins:
*         ___
*   1 o---UUU---o 2
*
*----------------------------------------------
* 
*  Equivalent circuit:
*
*         L1         R1
*    (1)  ___  (3)   ___  (2)
*     o-o-UUU---o---|___|-o-o
*       |                 |
*       |                 |
*       |       C1 ||     |
*       o----------||-----o
*       |          ||     |
*       |                 |
*       |    R2 ___       |
*       '------|___|------'
*
*
* L1 = inductance
* R1 = equivalent series resistance
* C1 = equivalent parallel capacitance
* R2 = equivalent parallel resistance
* 
*----------------------------------------------
*
.SUBCKT L_LINEAR 1 2 PARAMS: Inductance=10e-6 Rs=0.01 Cp=2e-12 Rp=300e3
*
L1 1 3 {Inductance}
R1 3 2 {Rs}
C1 1 2 {Cp}
R2 1 3 {Rp}
.ENDS L_LINEAR
