* This subcircuit line has no pins:
.SUBCKT shorty
.ends shorty