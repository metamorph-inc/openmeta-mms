*----------------------------------------------------------------------
* 2x8_header.cir
*
* SPICE Netlist: 8-pin header, 1x8, 2.54mm pitch, 5.08mm row spacing
*
* Copyright(C) 2014 MetaMorph Inc.
* http://metamorphsoftware.com/
*
*
*----------------------------------------------------------------------
* One row may be used as an 8-pin Arduino shield connector, the other
* row as corresponding test points.
*----------------------------------------------------------------------
*
*
*
*
*
*      (PIN1)  R1 ___
*         o------|___|----.
*                         |
*      (PIN2)  R2 ___     |
*         o------|___|----+
*                         |
*      (PIN3)  R3 ___     |
*         o------|___|----+
*                         |
*      (PIN4)  R4 ___     |
*         o------|___|----+
*                         |
*      (PIN5)  R5 ___     |
*         o------|___|----+
*                         |
*      (PIN6)  R6 ___     |
*         o------|___|----+
*                         |
*      (PIN7)  R7 ___     |
*         o------|___|----+
*                         |
*      (PIN8)  R8 ___     |
*         o------|___|----+
*                         |
*                         |
*                      (0)|
*                        ===
*                        GND
*
*
*
* PIN1 - PIN 8: -- External pins
*
* R1 - R8: -- 10^12 ohms; Leakage resistance of mounted pin to ground.
*
*
*----------------------------------------------------------------------
.SUBCKT HEADER_1X8 PIN1 PIN2 PIN3 PIN4 PIN5 PIN6 PIN7 PIN8
*
R1  PIN1 0    10E12
R2  PIN2 0    10E12
R3  PIN3 0    10E12
R4  PIN4 0    10E12
R5  PIN5 0    10E12
R6  PIN6 0    10E12
R7  PIN7 0    10E12
R8  PIN8 0    10E12
.ENDS 1X8_HEADER


