*----------------------------------------------------------------------
* res_0603.cir
*
* SPICE Netlist: Resistor chip, 0603 package
*
* Copyright(C) 2014 MetaMorph Inc.
* http://metamorphsoftware.com/
*
*
*----------------------------------------------------------------------
* This circuit is used to test SPICE model importing via CAT.
*----------------------------------------------------------------------
* 
* 
* 
*        (1)
*         o-----------.
*                     |
*                     | L1
*                     C|
*                     C|
*                     C|
*                     |
*                     | (11)
*                     |
*                     |
*                     | R1
*                    .-.
*                    | |
*                    | |
*                    '-'
*                     |
*        (2)          |
*         o-----------'
* 
* 
*   
*----------------------------------------------------------------------
.SUBCKT RES_0603 1 2 RVAL=1.0k
L1  1 11 800pH
R1 11  2 RVAL
.ENDS RES_0603


