RC time delay circuit
v1 1 0 dc 10
c1 1 2 47u ic=0
c2 1 2 22u ic=0
r1 2 3 3.3k
r2 3 4 3.3k
r3 4 5 3.3k
r4 5 6 3.3k
r5 6 7 3.3k
r6 7 8 3.3k
r7 8 9 3.3k
r8 9 10 3.3k
r9 10 11 3.3k
r10 11 12 3.3k
r11 12 13 3.3k
r12 13 14 3.3k
r13 14 15 3.3k
r14 15 16 3.3k
r15 16 17 3.3k
r16 17 18 3.3k
r17 18 19 3.3k
r18 19 20 3.3k
r19 20 21 3.3k
r20 21 22 3.3k
r21 22 23 3.3k
r22 23 24 3.3k
r23 24 25 3.3k
r24 25 26 3.3k
r25 26 27 3.3k
r26 27 28 3.3k
r27 28 29 3.3k
r28 29 30 3.3k
r29 30 31 3.3k
r30 31 32 3.3k
r31 32 33 3.3k
r32 33 34 3.3k
r33 34 35 3.3k
r34 35 36 3.3k
r35 36 37 3.3k
r36 37 38 3.3k
r37 38 39 3.3k
r38 39 40 3.3k
r39 40 41 3.3k
r40 41 42 3.3k
r41 42 43 3.3k
r42 43 44 3.3k
r43 44 45 3.3k
r44 45 46 3.3k
r45 46 47 3.3k
r46 47 48 3.3k
r47 48 49 3.3k
r48 49 50 3.3k
r49 50 0 3.3k
.tran 1nS 0.0032
.end 