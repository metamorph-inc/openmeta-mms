* INMP401 MEMS Microphone SPICE Model
.SUBCKT INMP401 VDD GND OUT
E1 N001 0 VDD GND 0.5
R1 N001 OUT 200
R2 VDD GND 13k
R3 OUT 0 18k
.ENDS INMP401