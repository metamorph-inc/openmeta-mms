*************************************************************
* Ngspice .cir file for C_TANT_0805_10u_10V_10%_AVX
*************************************************************
* AVX Tantalum Capacitor TAJP106K010R
*
.SUBCKT TAJP106K010R POS NEG

*PARASITIC INDUCTANCE
LESL POS 2 2.400000E-009
RELS POS 2 10

*LEAKAGE CURRENT & REVERSE BIAS EFFECTS
RP 2 NEG 1.100000E+007
DP NEG 2 DFWD

*RC-LADDER MODEL OF FREQUENCY EFFECTS
R1 2 3 RMOD1 2.881150E+000
C1 2 3 CMOD1 1.940236E-004
R2 3 4 RMOD2 9.540978E-001
C2 4 NEG CMOD2 3.242025E-007
R3 4 5 RMOD3 5.086542E-001
C3 5 NEG CMOD3 6.484049E-007
R4 5 6 RMOD4 2.541554E-001
C4 6 NEG CMOD4 1.296810E-006
R5 6 7 RMOD5 1.012703E+000
C5 7 NEG CMOD5 2.593620E-006
R6 7 8 RMOD6 4.602637E+000
C6 8 NEG CMOD6 5.187239E-006

.MODEL CMOD1 C (TNOM=25 TC1=1.463615E-003 TC2=-4.147800E-005)
.MODEL CMOD2 C (TNOM=25 TC1=3.749220E-004 TC2=2.806000E-006)
.MODEL CMOD3 C (TNOM=25 TC1=3.749220E-004 TC2=2.806000E-006)
.MODEL CMOD4 C (TNOM=25 TC1=3.749220E-004 TC2=2.806000E-006)
.MODEL CMOD5 C (TNOM=25 TC1=3.749220E-004 TC2=2.806000E-006)
.MODEL CMOD6 C (TNOM=25 TC1=3.749220E-004 TC2=2.806000E-006)
.MODEL RMOD1 R (TNOM=25 TC1=5.948893E-003 TC2=5.337100E-005)
.MODEL RMOD2 R (TNOM=25 TC1=-1.770874E-003 TC2=1.281300E-005)
.MODEL RMOD3 R (TNOM=25 TC1=-7.138201E-003 TC2=2.153200E-005)
.MODEL RMOD4 R (TNOM=25 TC1=-7.138201E-003 TC2=2.153200E-005)
.MODEL RMOD5 R (TNOM=25 TC1=-7.138201E-003 TC2=2.153200E-005)
.MODEL RMOD6 R (TNOM=25 TC1=-7.138201E-003 TC2=2.153200E-005)
.MODEL DFWD D (RS=0.1 IS=8E-10 N=2.5 XTI=0 EG=0.1)

.ENDS TAJP106K010R
*************************************************************
