* Hack for Connector Split
* connections:      Port B 0 .. B7
*                   |   
*                   |                        |   B0  .... B
*                   |   
.SUBCKT split8Bit      1   2   3 4 5 6 7 8   11 12 13 14 15 16 17 18 

R0 1 11 0.001
R1 2 12 0.001
R2 3 13 0.001
R3 4 14 0.001
R4 5 15 0.001
R5 6 16 0.001
R6 7 17 0.001
R7 8 18 0.001

.ENDS split8Bit
