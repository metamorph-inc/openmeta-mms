* NPN Transistor 2N2222 
* connections:      Collector
*                   |   Base
*                   |   |   Emitter
*                   |   |   |
.SUBCKT NPN2N222    1   2   3
Qxx 1 2 3 Q2N222A
.model Q2N222A NPN (IS=14.34F XTI=3 EG=1.11 VAF= 74.03 BF=255.9 NE=1.307 ISE=14.34F IKF=.2847 XTB=1.5 BR=6.092 NC=2 ISC=0 IKR=0 RC=1 CJC=7.306P MJC=.3416 VJC=.75 FC=.5 CJE=22.01P MJE=.377 VJE=.75 TR=46.91N TF=411.1P ITF=.6 VTF=1.7 XTF=3 RB=10) 
.ENDS NPN2N222
