* Lite-on LED

.MODEL D_green D (IS=575u  RS=25 N=6.79 BV=5 IBV=30U CJO=50P VJ=.75 M=150 )