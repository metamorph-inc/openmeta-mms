* R_CHIP
* Simple generic SPICE model of a chip resistor.
*
*
*----------------------------------------------
*  External Pins:
*
*   1 ---/\/\/\/\--- 2
*
*----------------------------------------------
* 
*  Equivalent circuit:
*
*                 C1
* 
*                 ||
*       .---------||--------.
*       |         ||        |
*       |   R1         L1   |
*   (1) |   ___   (3)  ___  | (2)
*     o-o--|___|---o---UUU--o-o
*
* R1 = "Resistance"
* L1 = "Ls"
* C1 = "Cp"
* 
*----------------------------------------------
*
.SUBCKT R_CHIP 1 2 PARAMS: Resistance=1k Ls=0.2e-12 Cp=280p
R1 1 3 {Resistance}
L1 3 2 {Ls}
C1 1 2 {Cp}
.ENDS R_CHIP